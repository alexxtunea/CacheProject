module fsm(
    input clk, rst, beg,
    input write,
    input read,
    input hit, miss,
    input free,
    output reg c0,c1,c2,c3,c4,c5,c6,c7
);

//FSM States 
parameter IDLE = 4'b0000;
parameter READ = 4'b0001;
parameter WRITE = 4'b0010;
parameter READ_HIT = 4'b0011;
parameter READ_MISS = 4'b0100;
parameter WRITE_HIT = 4'b0101;
parameter WRITE_MISS = 4'b0110;
parameter CHECK = 4'b0111;
parameter EVICT = 4'b1000;
parameter EXIT = 4'b1001;

reg [3:0] st, nxt_st;


always @(posedge clk,negedge rst) begin

    if(rst) begin
        st <= IDLE;
        {c0, c1, c2, c3, c4, c5, c6, c7} <= 8'b0;
    end
    else begin
        st <= nxt_st;
    end

end


always @(*) begin
    nxt_st = st;
    case(st)
        IDLE : begin
            if(bgn == 1'b0)begin
                nxt_state <= IDLE;
            end
            else begin
		if(read == 1'b1) begin
                nxt_st <= READ;
           	end
            	else if(write == 1'b1) begin
                nxt_st <= WRITE;
            	end
            	else begin
                nxt_st <= IDLE;
            	end
	    end     	
        end
        READ : begin
            if(hit == 1'b1) begin
                nxt_st <= READ_HIT;
            end
            else if(miss == 1'b1) begin
                nxt_st <= READ_MISS;
                
            end
        end
        WRITE : begin
            if(hit == 1'b1) begin
                nxt_st <= WRITE_HIT;
            end
            else if(miss == 1'b1) begin
                nxt_st <= WRITE_MISS;
            end
        end
        READ_HIT : begin
            nxt_st <= IDLE;
        end
        WRITE_HIT : begin
            nxt_st <= IDLE;
        end
        WRITE_MISS : begin
            nxt_st <= CHECK;
        end
        READ_MISS : begin
            nxt_st <= CHECK;
        end
        CHECK : begin 
            if(full == 1'b0) begin
                nxt_st <= EXIT;
            end
            if(full == 1'b1) begin
                nxt_st <= EVICT;
            end
        end
        EVICT : begin
            nxt_st <= EXIT;
        end
        EXIT : begin
            nxt_st <= IDLE;
        end

    endcase
end


always @(posedge clk,posedge rst) begin
    {c0, c1, c2, c3, c4, c5, c6, c7} <= 8'b0;

    case(nxt_st)
        IDLE : begin
            c0 <= 1'b1;
        end
        READ : begin
            c1 <= 1'b1;
        end
        WRITE : begin
            c2 <= 1'b1;
        end
        READ_HIT : begin
            c1 <= 1'b1;
            c3 <= 1'b1;
        end
        WRITE_HIT : begin
            c2 <= 1'b1;
            c3 <= 1'b1;
        end
        READ_MISS : begin
            c1 <= 1'b1;
            c4 <= 1'b1;
        end
        WRITE_MISS : begin
            c2 <= 1'b1;
            c4 <= 1'b1;
        end
        CHECK : begin
            c5 <= 1'b1;
        end
        EVICT : begin
            c7 <= 1'b1;
        end
        EXIT : begin
            c6 <= 1'b1;
        end
    endcase
end

endmodule


module Cache #(
     parameter CACHE_SIZE = 32768, //32 KB
     parameter BLOCK_SIZE = 64, //64 bytes for each block
     parameter NO_SETS = 128, //numarul de seturi 
     parameter CACHE_TYPE = 4, // 4 way associativity
     parameter WORD_SIZE = 4 //each word has 4 bytes 
)(
     input clk, rst,
     input c0,c1,c2,c3,c4,c5,c6,c7,
     input [31:0] address, 
     input [511:0] data_to_write,
     input read, write,
     output reg [511:0] read_data,
     output reg [3:0] dirty,
     output reg [3:0] and_val,
     output reg hit, miss, free
);

parameter NO_BLOCKS = BLOCK_SIZE / WORD_SIZE;
parameter INDEX_BITS = $clog2(NO_SETS);
parameter OFFSET_BITS = $clog2(BLOCK_SIZE);
parameter TAG_BITS = 32 - (INDEX_BITS + OFFSET_BITS);


reg [NO_SETS*CACHE_TYPE-1:0] data_cache[NO_SETS*CACHE_TYPE-1:0];
reg [TAG_BITS-1:0] tags_cache[NO_SETS*CACHE_TYPE-1:0];
reg [NO_SETS*CACHE_TYPE-1:0] valid;
reg [CACHE_TYPE-1:0] dirty_bits[NO_SETS*CACHE_TYPE-1:0];
reg [CACHE_TYPE + $clog2(CACHE_TYPE) -1 :0] lru[NO_SETS-1:0];

reg [INDEX_BITS- 1:0] index;
reg [OFFSET_BITS-1:0] offset;
reg [TAG_BITS-1:0] tag;
integer i, j, way_set, br;


//temporary values 
reg [511:0] data_from_cache;
reg [3:0] temp_tag;
reg [3:0] temp_and_values;
reg temp_hit;
reg [1:0] pos_for_new_data;

reg [1:0] st, st_next;

    always @(posedge clk,negedge rst) begin
        if(c0 == 1'b1) begin
            tag <= address[31:13];
            index <= address[12:6];
            offset <= address[5:0];
            
        end
    end

 always @(posedge clk,negedge rst) begin

        if(tag == tags_cache[index]) begin
            temp_tag[0] <= 1'b1;
        end
        else begin
            temp_tag[0] <= 1'b0;
        end
        //tag for set 3
        if(tag == tags_cache[128+index]) begin
            temp_tag[1] <= 1'b1;
        end
        else begin
            temp_tag[1] <= 1'b0;
        end
        //tag for set 2
        if(tag == tags_cache[2*128+index]) begin
            temp_tag[2] <= 1'b1;
        end
        else begin
            temp_tag[2] <= 1'b0;
        end
        //tag for set 1
        if(tag == tags_cache[3*128+index]) begin
            
            temp_tag[3] <= 1'b1;
        end
        else begin
            temp_tag[3] <= 1'b0;
        end

        //AND operations between comparator and valid
        temp_and_values[3] <= temp_tag[3] && valid[3*128+index];
        temp_and_values[2] <= temp_tag[2] && valid[2*128+index];
        temp_and_values[1] <= temp_tag[1] && valid[128+index];
        temp_and_values[0] <= temp_tag[0] && valid[index];

         
        //OR operation between AND gates
        temp_hit <= temp_and_values[0] || temp_and_values[1] || temp_and_values[2] || temp_and_values[3];


        //MUX 4:1
        if(temp_and_values[3] == 1'b1) begin
            data_from_cache <= data_cache[3*128+index][511:0];
        end
        if(temp_and_values[2] == 1'b1) begin
            data_from_cache <= data_cache[2*128+index][511:0];
            
        end
        if(temp_and_values[1] == 1'b1) begin
            data_from_cache <= data_cache[128+index][511:0];
            
        end
        if(temp_and_values[0] == 1'b1) begin
            data_from_cache <= data_cache[index][511:0]; 
        end
        
    end

always @(posedge clk,negedge rst) begin
        hit <= 1'b0;
	miss <= 1'b0;

        if(rst) begin

            valid <= 512'b0;

            for (i = 0; i < 128; i = i + 1) begin
                lru[i] <= 12'b100100100100;
                   
            end
        end
        else begin
            if(st == ) begin //read


                if(temp_hit == 4'b0) begin
                    hit <= 1'b0;
		    miss <= 1'b1;
                end
                else begin
                    hit <= 1'b0;
		    miss <= 1'b1;		    

                    //for dirty bit when you get the second hit from the same data
                    //set1
                    if(temp_and_values[3] == 1'b1 && dirty_bits[index][3] == 1'b0) begin
                        dirty_bits[index][3] <= 1'b1;
                    end
                    //set2
                    if(temp_and_values[2] == 1'b1 && dirty_bits[index][2] == 1'b0) begin
                        dirty_bits[index][2] <= 1'b1;               
                    end
                    //set3
                    if(temp_and_values[1] == 1'b1 && dirty_bits[index][1] == 1'b0) begin
                        dirty_bits[index][1] <= 1'b1;
                    end
                    //set4
                    if(temp_and_values[0] == 1'b1 && dirty_bits[index][0] == 1'b0) begin
                        dirty_bits[index][0] <= 1'b1;
                    end
                end

                dirty <= dirty_bits[index];

                if(c3 == 1'b1) begin
                    outbus <= data_from_cache;
                end

                and_val <= temp_and_values; // shows in which set was stored data
            end
            if(c2 == 1'b1) begin //write
         
                if(temp_hit == 4'b0) begin
                    hit <= 1'b0;
		    miss <= 1'b1;
                end
                else begin
                    hit <= 1'b0;
		    miss <= 1'b1;

                    //for dirty bit when you get the second hit from the same data 
                    //and when you need to send data to the main memory
                    //set1
                    if(temp_and_values[3] == 1'b1 && dirty_bits[index][3] == 1'b0 && c3 == 1'b1) begin
                        dirty_bits[index][3] <= 1'b1;
                        read_data <= data_from_cache;
                    end
                    //set2
                    if(temp_and_values[2] == 1'b1 && dirty_bits[index][2] == 1'b0 && c3 == 1'b1) begin
                        dirty_bits[index][2] <= 1'b1;
                        read_data <= data_from_cache;               
                    end
                    //set3
                    if(temp_and_values[1] == 1'b1 && dirty_bits[index][1] == 1'b0 && c3 == 1'b1) begin
                        dirty_bits[index][1] <= 1'b1;
                        read_data <= data_from_cache;
                    end
                    //set4
                    if(temp_and_values[0] == 1'b1 && dirty_bits[index][0] == 1'b0 && c3 == 1'b1) begin
                        dirty_bits[index][0] <= 1'b1;
                        read_data <= data_from_cache;
                    end
                    dirty <= dirty_bits[index];
                end

                and_val <= temp_and_values;// shows in which set was stored data
                
            end
            if(c6 == 1'b1) begin //Load the date into the cache
                

                if(pos_for_new_data == 2'b11) begin
                    lru[index][11:9] <= 3'b000;
                    dirty_bits[index][3] <= 1'b0;
                    data_cache[3*128+index] <= data;
                    tags_cache[3*128+index] <= tag;
                    valid[3*128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b10) begin
                    lru[index][8:6] <= 3'b000;
                    dirty_bits[index][2] <= 1'b0;
                    data_cache[2*128+index] <= data;
                    tags_cache[2*128+index] <= tag;
                    valid[2*128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b01) begin
                    lru[index][5:3] <= 3'b000;
                    dirty_bits[index][1] <= 1'b0;
                    data_cache[128+index] <= data;
                    tags_cache[128+index] <= tag;
                    valid[128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b00) begin
                    lru[index][2:0] <= 3'b000;
                    dirty_bits[index][0] <= 1'b0;
                    data_cache[index] <= data;
                    tags_cache[index] <= tag;
                    valid[index] <= 1'b1;
                end
                
            end

        end
    end

	
endmodule




















