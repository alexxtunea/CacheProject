'import "fsm.v"

module Cache #(
     parameter CACHE_SIZE = 32768, //32 KB
     parameter BLOCK_SIZE = 64, //64 bytes for each block
     parameter NO_SETS = 128, //numarul de seturi 
     parameter CACHE_TYPE = 4, // 4 way associativity
     parameter WORD_SIZE = 4 //each word has 4 bytes 
)(
     input clk, rst,
     input c0,c1,c2,c3,c4,c5,c6,c7,
     input [31:0] address, 
     input [511:0] data_to_write,
     input read, write, 
     output reg [511:0] read_data,
     output reg [3:0] dirty,
     output reg [3:0] and_val,
     output reg hit, miss, free, ask_for_data
);

parameter NO_BLOCKS = BLOCK_SIZE / WORD_SIZE;
parameter INDEX_BITS = $clog2(NO_SETS);
parameter OFFSET_BITS = $clog2(BLOCK_SIZE);
parameter TAG_BITS = 32 - (INDEX_BITS + OFFSET_BITS);


reg [NO_SETS*CACHE_TYPE-1:0] data_cache[NO_SETS*CACHE_TYPE-1:0];
reg [TAG_BITS-1:0] tags_cache[NO_SETS*CACHE_TYPE-1:0];
reg [NO_SETS*CACHE_TYPE-1:0] valid;
reg [CACHE_TYPE-1:0] dirty_bits[NO_SETS*CACHE_TYPE-1:0];
reg [CACHE_TYPE + $clog2(CACHE_TYPE) -1 :0] lru[NO_SETS-1:0];

reg [INDEX_BITS- 1:0] index;
reg [OFFSET_BITS-1:0] offset;
reg [TAG_BITS-1:0] tag;
integer i, j, way_set, br;


//temporary values 
reg [511:0] data_from_cache;
reg [3:0] temp_tag;
reg [3:0] temp_and_values;
reg temp_hit;
reg [1:0] new_location;

reg [1:0] st, st_next;

    always @(posedge clk,negedge rst) begin
        if(c0 == 1'b1) begin
            tag <= address[31:13];
            index <= address[12:6];
            offset <= address[5:0];
            
        end
    end

 always @(posedge clk,negedge rst) begin

	   for(i=0; i < CACHE_TYPE; i = i + 1) begin: gen_temp_tag
		if(tag == tags_cache[NO_SETS * i + index]) begin
			temp_tag[i] <= 1'b1;
		end
		else begin
			temp_tag[i] <= 1'b0;
		end
           end


	   for(i=CACHE_TYPE-1; i>=0; i = i-1) begin: gen_tempvalues_temphit
		temp_and_values[i] <= temp_tag[i] && valid[i*NO_SETS+index];
		temp_hit <= temp_hit || temp_and_values[i];
	   end
         
	
        //MUX 4:1
	   for(i = CACHE_TYPE - 1; i >= 0; i = i - 1) begin: gen_tempvalues
		if(temp_and_values[i] == 1'b1) begin
		   data_from_cache <= data_cache[i*NO_SETS+index][NO_SETS*CACHE_TYPE-1:0];
		end
	   end
                
end

always @(posedge clk,negedge rst) begin
        hit <= 1'b0;
	miss <= 1'b0;

        if(rst) begin

            valid <= 512'b0;

            for (i = 0; i < NO_SETS; i = i + 1) begin
                lru[i] <= 12'b100100100100;
                   
            end
        end
        else begin
            if(c1 == 1'b1) begin //read
                if(temp_hit == 4'b0) begin
                    hit <= 1'b0;
		    miss <= 1'b1;
                end
                else begin
                    hit <= 1'b0;
		    miss <= 1'b1;		    

                    //for dirty bit when you get the second hit from the same data
			for(i = CACHE_TYPE - 1; i>=0; i = i-1) begin
				if(temp_and_values[i] == 1'b1 && dirty_bits[index][i] == 1'b0) begin
                        		dirty_bits[index][i] <= 1'b1;
				end
			end
                end

                dirty <= dirty_bits[index];

                if(c3 == 1'b1) begin
                    read_data <= data_from_cache;
                end

                and_val <= temp_and_values; // shows in which set was stored data
            end
            if(c2 == 1'b1) begin //write
         
                if(temp_hit == 4'b0) begin
                    hit <= 1'b0;
		    miss <= 1'b1;
                end
                else begin
                    hit <= 1'b0;
		    miss <= 1'b1;

                    //for dirty bit when you get the second hit from the same data 
                    //and when you need to send data to the main memory
                    //set1

		
		    for(i = CACHE_TYPE - 1; i >= 0; i = i-1) begin
			if(temp_and_values[i] == 1'b1 && dirty_bits[index][i] == 1'b0 && c3 == 1'b1) begin
                        	dirty_bits[index][i] <= 1'b1;
                        	read_data <= data_from_cache;
                    	end
		    end
                    
                    dirty <= dirty_bits[index];
                end

                and_val <= temp_and_values;// shows in which set was stored data
                
            end
            if(c6 == 1'b1) begin //Load the date into the cache
                
                if(pos_for_new_data == 2'b11) begin
                    lru[index][11:9] <= 3'b000;
                    dirty_bits[index][3] <= 1'b0;
                    data_cache[3*128+index] <= data_to_write;
                    tags_cache[3*128+index] <= tag;
                    valid[3*128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b10) begin
                    lru[index][8:6] <= 3'b000;
                    dirty_bits[index][2] <= 1'b0;
                    data_cache[2*128+index] <= data_to_write;
                    tags_cache[2*128+index] <= tag;
                    valid[2*128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b01) begin
                    lru[index][5:3] <= 3'b000;
                    dirty_bits[index][1] <= 1'b0;
                    data_cache[128+index] <= data_to_write;
                    tags_cache[128+index] <= tag;
                    valid[128+index] <= 1'b1;
                end
                else if(pos_for_new_data == 2'b00) begin
                    lru[index][2:0] <= 3'b000;
                    dirty_bits[index][0] <= 1'b0;
                    data_cache[index] <= data_to_write;
                    tags_cache[index] <= tag;
                    valid[index] <= 1'b1;
                end
                
            end

        end
    end

    always @(posedge clk, negedge rst) begin
	if(c4 == 1'b1) begin
		ask_for_data <= 1'b1;
	end
	else begin
            ask_for_data <= 1'b0;
        end
    end

    //LRU
    always @(posedge clk,negedge rst) begin
        if(c3 == 1'b1) begin
            //When you get a hit and reset the LRU data to 0 and increment the over LRU data
            if(temp_and_values == 4'b1000) begin //set1
                lru[index][11:9] <= 3'b0;
                if(lru[index][8:6] < 3'b011) begin
                    lru[index][8:6] <= lru[index][8:6] + 3'b001;
                end
                if(lru[index][5:3] < 3'b011) begin
                    lru[index][5:3] <= lru[index][5:3] + 3'b001;
                end
                if(lru[index][2:0] < 3'b011) begin
                    lru[index][2:0] <= lru[index][2:0] + 3'b001;
                end

            end 
            else if(temp_and_values == 4'b0100) begin //set2
                lru[index][8:6] <= 3'b0;
                if(lru[index][11:9] < 3'b011) begin
                    lru[index][11:9] <= lru[index][11:9] + 3'b001;
                end
                if(lru[index][5:3] < 3'b011) begin
                    lru[index][5:3] <= lru[index][5:3] + 3'b001;
                end
                if(lru[index][2:0] < 3'b011) begin
                    lru[index][2:0] <= lru[index][2:0] + 3'b001;
                end
            end
            else if(temp_and_values == 4'b0010) begin //set3
                lru[index][5:3] <= 3'b0;
                if(lru[index][8:6] < 3'b011) begin
                    lru[index][8:6] <= lru[index][8:6] + 3'b001;
                end
                if(lru[index][11:9] < 3'b011) begin
                    lru[index][11:9] <= lru[index][11:9] + 3'b001;
                end
                if(lru[index][2:0] < 3'b011) begin
                    lru[index][2:0] <= lru[index][2:0] + 3'b001;
                end
            end
            else if(temp_and_values == 4'b0001) begin //set4
                lru[index][2:0] <= 3'b0;
                if(lru[index][8:6] < 3'b011) begin
                    lru[index][8:6] <= lru[index][8:6] + 3'b001;
                end
                if(lru[index][5:3] < 3'b011) begin
                    lru[index][5:3] <= lru[index][5:3] + 3'b001;
                end
                if(lru[index][11:9] < 3'b011) begin
                    lru[index][11:9] <= lru[index][11:9] + 3'b001;
                end
            end
        end

        if(c5 == 1'b1) begin
            
            //When you get a miss and need to give a position for the next data if there
            //is space in cache
            if(lru[index][11:9] == 3'b100) begin
                new_location <= 2'b11;
                space_in_lru <= 1'b0;
                
            end
            else if(lru[index][8:6] == 3'b100) begin
                new_location <= 2'b10;
                space_in_lru <= 1'b0;
                
            end
            else if(lru[index][5:3] == 3'b100) begin
                new_location <= 2'b01;
                space_in_lru <= 1'b0;
                
            end
            else if(lru[index][2:0] == 3'b100) begin
                new_location <= 2'b00;
                space_in_lru <= 1'b0;
                
            end
            else begin
                space_in_lru <= 1'b1;
                
            end
            
        end

        if(c7 == 1'b1) begin
            //makes space in cache when everything is full by giving the position 
            //of the last reacent used set
            if(lru[index][11:9] == 3'b011) begin
                new_location <= 2'b11;
            end
            else if(lru[index][8:6] == 3'b011) begin
                new_location <= 2'b10;
            end
            else if(lru[index][5:3] == 3'b011) begin
                new_location <= 2'b01;
            end
            else if(lru[index][2:0] == 3'b011) begin
                new_location <= 2'b00;
            end
            
        end 
        
    end

	
endmodule




















